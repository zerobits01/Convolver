library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity non_pipeline_convolver is
end non_pipeline_convolver;

architecture Behavioral of non_pipeline_convolver is

begin


end Behavioral;

