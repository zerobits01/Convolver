library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library work;
use work.arr_mat.all;

entity PAM_TOP is
	Port(
		
	);
end PAM_TOP;

architecture Behavioral of PAM_TOP is

begin


end Behavioral;

