library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Arr_Mat is

	type int_arr is array(0 to 90) of integer;
	type int_mat is array(0 to 10) of int_arr;
end Arr_Mat;

package body Arr_Mat is

end Arr_Mat;
